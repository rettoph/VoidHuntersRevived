entity:ship-part:hull:hexagonentity:ship-part:hull:square  entity:ship-part:hull:triangle entity:ship-part:hull:square  entity:ship-part:hull:hexagon  entity:ship-part:hull:square  entity:ship-part:hull:triangle entity:ship-part:hull:square   #entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driverentity:ship-part:hull:square #entity:ship-part:weapon:mass-driver     entity:ship-part:hull:square  entity:ship-part:hull:triangle entity:ship-part:hull:square  entity:ship-part:hull:hexagon  entity:ship-part:hull:square  entity:ship-part:hull:triangle  #entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver    entity:ship-part:hull:square  entity:ship-part:hull:triangle entity:ship-part:hull:square  entity:ship-part:hull:hexagon  entity:ship-part:hull:square  entity:ship-part:hull:triangle entity:ship-part:hull:square   #entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver    entity:ship-part:hull:square  entity:ship-part:hull:triangle entity:ship-part:hull:square  entity:ship-part:hull:hexagon  entity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:hull:triangle entity:ship-part:hull:square entity:ship-part:thruster:small entity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:small#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver    entity:ship-part:hull:square  entity:ship-part:hull:triangle entity:ship-part:hull:square  entity:ship-part:hull:hexagon  entity:ship-part:hull:square  entity:ship-part:hull:triangle entity:ship-part:hull:square   #entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver    entity:ship-part:hull:square  entity:ship-part:hull:triangle entity:ship-part:hull:square  entity:ship-part:hull:hexagon  entity:ship-part:hull:square  entity:ship-part:hull:triangle entity:ship-part:hull:square   #entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver    