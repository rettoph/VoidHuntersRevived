 Unnamed Ship!entity:ship-part:chassis:mosquito  entity:ship-part:thruster:smallentity:ship-part:thruster:small    entity:ship-part:thruster:small  