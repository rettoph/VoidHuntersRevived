 Unnamed Shipchassis:mosquitothruster:smallthruster:smallthruster:smallthruster:smallthruster:smallthruster:small hull:pentagon   weapon:gun:mass-driver weapon:gun:mass-driverhull:pentagon  weapon:gun:mass-driver   