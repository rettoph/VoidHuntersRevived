ship-part:hexagonship-part:pentagon  ship-part:square  ship-part:hexagon  ship-part:square  ship-part:triangle  ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:square ship-part:weapon:mass-driver     ship-part:pentagon  ship-part:square  ship-part:hexagon  ship-part:square  ship-part:triangle  ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:square ship-part:weapon:mass-driver     ship-part:pentagon  ship-part:square  ship-part:hexagon  ship-part:square  ship-part:triangle  ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:square ship-part:weapon:mass-driver     ship-part:pentagon  ship-part:square  ship-part:hexagon  ship-part:square  ship-part:triangle  ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:square ship-part:weapon:mass-driver     ship-part:pentagon  ship-part:square  ship-part:hexagon  ship-part:square  ship-part:triangle  ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:square ship-part:weapon:mass-driver     ship-part:pentagon  ship-part:square  ship-part:hexagon  ship-part:square  ship-part:triangleship-part:weapon:mass-driver ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:square ship-part:weapon:mass-driver     ship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:weapon:mass-drivership-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:squareship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:squareship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:squareship-part:thruster:smallship-part:squareship-part:thruster:smallship-part:squareship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:squareship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:weapon:mass-drivership-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:squareship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:squareship-part:thruster:smallship-part:squareship-part:thruster:smallship-part:squareship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:squareship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:weapon:mass-drivership-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:pentagonship-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:thruster:smallship-part:pentagonship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:thruster:smallship-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:smallship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:squareship-part:weapon:mass-drivership-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:squareship-part:weapon:mass-drivership-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:thruster:smallship-part:pentagonship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:thruster:smallship-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:smallship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:squareship-part:weapon:mass-drivership-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:squareship-part:weapon:mass-drivership-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-driver ship-part:thruster:small