 Unnamed Shipvhr:chassis:squid vhr:hull:square vhr:weapon:mass-driver  vhr:weapon:mass-drivervhr:weapon:mass-driver vhr:hull:square vhr:weapon:mass-driver     vhr:thruster:smallvhr:thruster:small  vhr:thruster:smallvhr:thruster:small