 Unnamed Shipvhr:chassis:bullfrogvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:thruster:small vhr:hull:lattice vhr:weapon:mass-driver     vhr:thruster:small vhr:thruster:smallvhr:thruster:small vhr:weapon:mass-drivervhr:weapon:mass-drivervhr:hull:lattice vhr:thruster:small     vhr:weapon:mass-driver vhr:thruster:smallvhr:thruster:small