 Unnamed Shipvhr:chassis:fightervhr:weapon:laser:tinyvhr:thruster:tinyvhr:thruster:tinyvhr:thruster:tinyvhr:thruster:tiny