 Unnamed Shipchassis:pelicanhull:diamond    thruster:small   armor:shield hull:diamond  thruster:small      thruster:smallweapon:gun:mass-driverweapon:gun:mass-driver armor:shield weapon:gun:mass-driverweapon:gun:mass-driverthruster:small