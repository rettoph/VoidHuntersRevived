entity:ship-part:hull:triangleentity:ship-part:hull:square  entity:ship-part:hull:square entity:ship-part:hull:square  entity:ship-part:hull:triangle  #entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driverentity:ship-part:hull:square #entity:ship-part:weapon:mass-driverentity:ship-part:hull:triangle #entity:ship-part:weapon:mass-driver   entity:ship-part:hull:square  entity:ship-part:hull:square entity:ship-part:hull:square  entity:ship-part:hull:triangle  #entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driverentity:ship-part:hull:square #entity:ship-part:weapon:mass-driverentity:ship-part:hull:triangle #entity:ship-part:weapon:mass-driver   entity:ship-part:hull:square  entity:ship-part:hull:square entity:ship-part:hull:square  entity:ship-part:hull:triangle  #entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driverentity:ship-part:hull:square #entity:ship-part:weapon:mass-driverentity:ship-part:hull:triangle #entity:ship-part:weapon:mass-driver   