 Unnamed Shipvhr:chassis:butterflyvhr:thruster:smallvhr:thruster:small vhr:hull:beam:vertical  vhr:weapon:mass-driver vhr:thruster:smallvhr:thruster:smallvhr:thruster:small vhr:hull:beam:verticalvhr:special:power-cell       vhr:hull:beam:vertical vhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:weapon:mass-driver   vhr:thruster:small