 Unnamed Shipvhr:chassis:waspvhr:special:power-cellvhr:thruster:smallvhr:hull:beam:verticalvhr:hull:squarevhr:thruster:smallvhr:hull:beam:horizontalvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:special:power-cellvhr:thruster:small  vhr:thruster:smallvhr:thruster:smallvhr:special:power-cellvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:thruster:small  vhr:special:power-cell vhr:hull:beam:verticalvhr:thruster:small vhr:hull:beam:verticalvhr:hull:square vhr:hull:beam:horizontalvhr:weapon:laservhr:weapon:laservhr:weapon:laservhr:hull:square vhr:hull:square  vhr:weapon:laservhr:weapon:laservhr:special:power-cellvhr:thruster:smallvhr:thruster:smallvhr:thruster:small   vhr:thruster:smallvhr:thruster:smallvhr:thruster:small vhr:thruster:smallvhr:thruster:smallvhr:thruster:small vhr:special:shield-generatorvhr:special:shield-generatorvhr:special:shield-generatorvhr:thruster:small vhr:thruster:smallvhr:special:power-cell  vhr:special:shield-generatorvhr:special:shield-generatorvhr:hull:beam:verticalvhr:hull:squarevhr:thruster:smallvhr:hull:beam:horizontalvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:special:power-cell  vhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:special:power-cellvhr:thruster:smallvhr:thruster:smallvhr:special:power-cellvhr:special:shield-generator vhr:hull:beam:verticalvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:hull:beam:verticalvhr:hull:squarevhr:thruster:smallvhr:hull:beam:horizontalvhr:weapon:laservhr:weapon:laservhr:weapon:laservhr:special:power-cellvhr:hull:squarevhr:weapon:laser  vhr:thruster:smallvhr:thruster:small vhr:thruster:smallvhr:thruster:smallvhr:thruster:small      