 Unnamed Shipvhr:chassis:squidvhr:special:fighter-bay  vhr:weapon:mass-drivervhr:weapon:mass-driver      vhr:thruster:smallvhr:thruster:smallvhr:hull:square vhr:weapon:mass-driver vhr:hull:square vhr:weapon:mass-driver vhr:thruster:smallvhr:thruster:small