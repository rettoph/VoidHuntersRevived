 Unnamed Shipvhr:chassis:dragonfly   vhr:thruster:small vhr:thruster:small     vhr:weapon:mass-drivervhr:thruster:smallvhr:thruster:smallvhr:hull:wing:right  vhr:hull:triangle vhr:weapon:mass-driver vhr:thruster:small  vhr:hull:wing:left vhr:thruster:small vhr:hull:trianglevhr:weapon:mass-driver     