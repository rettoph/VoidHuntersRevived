ship-part:chassis:mosquitoship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:small ship-part:pentagonship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:small  ship-part:weapon:mass-drivership-part:triangle  ship-part:weapon:mass-drivership-part:pentagon ship-part:weapon:mass-driver ship-part:thruster:small part:pentagon  ship-part:thruster:smallship-part:thruster:smallship-part:thruster:small ip-part:thruster:small 