 Unnamed Shipvhr:chassis:butterflyvhr:thruster:smallvhr:thruster:smallvhr:special:shield-generator     vhr:special:shield-generatorvhr:thruster:small