 Unnamed Shipvhr:chassis:pelicanvhr:armor:shield vhr:thruster:small vhr:thruster:smallvhr:weapon:mass-drivervhr:weapon:mass-driver vhr:armor:shield vhr:weapon:mass-drivervhr:weapon:mass-drivervhr:thruster:small vhr:thruster:small 