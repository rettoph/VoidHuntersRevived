 Unnamed Shipvhr:chassis:dragonflyvhr:thruster:smallvhr:thruster:smallvhr:special:power-cellvhr:special:power-cellvhr:thruster:smallvhr:special:power-cellvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:special:power-cellvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:hull:wing:right  vhr:hull:squarevhr:thruster:smallvhr:hull:wing:right  vhr:hull:wing:rightvhr:thruster:smallvhr:thruster:smallvhr:hull:trianglevhr:weapon:mass-drivervhr:hull:trianglevhr:hull:trianglevhr:weapon:mass-drivervhr:hull:trianglevhr:hull:trianglevhr:weapon:mass-drivervhr:thruster:small vhr:thruster:smallvhr:weapon:mass-drivervhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:special:power-cellvhr:thruster:smallvhr:thruster:smallvhr:hull:latticevhr:hull:latticevhr:hull:latticevhr:hull:latticevhr:hull:latticevhr:hull:latticevhr:hull:latticevhr:hull:latticevhr:hull:latticevhr:hull:latticevhr:hull:beam:horizontalvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:hull:triangle vhr:hull:trianglevhr:hull:squarevhr:special:power-cell vhr:thruster:smallvhr:thruster:smallvhr:thruster:small   vhr:special:fighter-bay   vhr:special:fighter-bay  vhr:special:fighter-bay   vhr:special:fighter-bay  vhr:hull:trianglevhr:special:shield-generatorvhr:thruster:smallvhr:thruster:small  vhr:special:fighter-bay  vhr:hull:triangle vhr:thruster:small   vhr:special:fighter-bay  vhr:special:fighter-bay   vhr:special:fighter-bay  vhr:special:fighter-bay   vhr:special:fighter-bay  vhr:special:fighter-bay   vhr:special:fighter-bay  vhr:special:fighter-bayvhr:thruster:small  vhr:special:fighter-bay  vhr:hull:triangle vhr:thruster:smallvhr:thruster:small  vhr:special:fighter-bay  vhr:hull:trianglevhr:special:shield-generatorvhr:thruster:small   vhr:special:fighter-bay vhr:thruster:smallvhr:hull:wing:leftvhr:hull:latticevhr:hull:latticevhr:hull:latticevhr:hull:latticevhr:hull:latticevhr:hull:latticevhr:hull:latticevhr:hull:latticevhr:hull:latticevhr:hull:latticevhr:hull:beam:horizontalvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:hull:trianglevhr:hull:trianglevhr:thruster:small     vhr:special:fighter-bay   vhr:special:fighter-bay  vhr:special:fighter-bay  vhr:thruster:smallvhr:special:fighter-bay  vhr:special:fighter-bay   vhr:hull:trianglevhr:thruster:smallvhr:special:shield-generator  vhr:special:fighter-bay   vhr:hull:trianglevhr:thruster:smallvhr:hull:beam:vertical vhr:special:shield-generatorvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:special:power-cellvhr:thruster:small  vhr:special:fighter-bay   vhr:special:fighter-bay  vhr:special:fighter-bay   vhr:special:fighter-bay  vhr:special:fighter-bay   vhr:special:fighter-bay  vhr:special:fighter-bay  vhr:thruster:smallvhr:special:fighter-bay  vhr:special:fighter-bay  vhr:thruster:smallvhr:hull:trianglevhr:thruster:smallvhr:hull:beam:vertical vhr:special:power-cellvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:special:shield-generatorvhr:thruster:small  vhr:special:fighter-bay   vhr:hull:trianglevhr:thruster:smallvhr:special:shield-generator vhr:thruster:smallvhr:thruster:smallvhr:hull:squarevhr:special:power-cellvhr:hull:wing:leftvhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:hull:wing:leftvhr:thruster:smallvhr:thruster:smallvhr:weapon:mass-drivervhr:hull:trianglevhr:hull:trianglevhr:thruster:smallvhr:hull:trianglevhr:hull:triangle vhr:hull:trianglevhr:thruster:smallvhr:weapon:mass-drivervhr:weapon:mass-drivervhr:weapon:mass-drivervhr:thruster:smallvhr:thruster:small  vhr:thruster:small  vhr:thruster:smallvhr:thruster:small