 Untitled Ship!entity:ship-part:chassis:mosquitoentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:small entity:ship-part:hull:pentagon  #entity:ship-part:weapon:mass-driver #entity:ship-part:weapon:mass-driverentity:ship-part:hull:pentagon #entity:ship-part:weapon:mass-driver   