 Unnamed Shipvhr:chassis:mosquitovhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:thruster:small vhr:hull:pentagon vhr:weapon:mass-driver  vhr:weapon:mass-drivervhr:hull:pentagon   vhr:weapon:mass-driver vhr:thruster:smallvhr:thruster:small