!entity:ship-part:chassis:mosquitoentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:small entity:ship-part:hull:pentagon  #entity:ship-part:weapon:mass-driver #entity:ship-part:weapon:mass-driverentity:ship-part:hull:pentagon #entity:ship-part:weapon:mass-driver   ship-part:hull:triangle     tity:ship-part:weapon:mass-driver   ity:ship-part:hull:square #entity:ship-part:weapon:mass-driverentity:ship-part:hull:triangle #entity:ship-part:weapon:mass-driverentity:ship-part:thruster:smallentity:ship-part:thruster:small entity:ship-part:hull:square  entity:ship-part:thruster:small  ip-part:weapon:mass-driver#entity:ship-part:weapon:mass-driverentity:ship-part:hull:square #entity:ship-part:weapon:mass-driverentity:ship-part:hull:triangle #entity:ship-part:weapon:mass-driverentity:ship-part:thruster:smallentity:ship-part:thruster:small :weapon:mass-driver#entity:ship-part:weapon:mass-driverentity:ship-part:hull:square #entity:ship-part:weapon:mass-driverentity:ship-part:hull:triangle #entity:ship-part:weapon:mass-driverentity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:hull:triangle entity:ship-part:hull:triangle #entity:ship-part:weapon:mass-driver entity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:small le entity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:thruster:small#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driverentity:ship-part:thruster:smallentity:ship-part:hull:square  entity:ship-part:hull:square entity:ship-part:hull:triangle entity:ship-part:thruster:smallentity:ship-part:hull:hexagon entity:ship-part:thruster:small entity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:hull:hexagon entity:ship-part:thruster:small entity:ship-part:hull:square entity:ship-part:hull:triangle entity:ship-part:thruster:small  #entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver  #entity:ship-part:weapon:mass-driver #entity:ship-part:weapon:mass-driverentity:ship-part:hull:triangle entity:ship-part:hull:hexagon  #entity:ship-part:weapon:mass-driverentity:ship-part:hull:square  entity:ship-part:hull:hexagon  #entity:ship-part:weapon:mass-driverentity:ship-part:hull:square #entity:ship-part:weapon:mass-driver entity:ship-part:hull:triangle  entity:ship-part:thruster:small entity:ship-part:thruster:smallentity:ship-part:thruster:small entity:ship-part:thruster:smallentity:ship-part:thruster:small entity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:hull:triangle #entity:ship-part:weapon:mass-driverentity:ship-part:hull:square #entity:ship-part:weapon:mass-driverentity:ship-part:thruster:smallentity:ship-part:thruster:small  -part:weapon:mass-driverentity:ship-part:hull:square #entity:ship-part:weapon:mass-driverentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:small entity:ship-part:weapon:mass-driver  #entity:ship-part:weapon:mass-driver #entity:ship-part:weapon:mass-driverentity:ship-part:hull:triangle entity:ship-part:hull:hexagon  #entity:ship-part:weapon:mass-driverentity:ship-part:hull:square  entity:ship-part:hull:hexagon  #entity:ship-part:weapon:mass-driverentity:ship-part:hull:square #entity:ship-part:weapon:mass-driver entity:ship-part:hull:triangle  entity:ship-part:thruster:small entity:ship-part:thruster:smallentity:ship-part:thruster:small entity:ship-part:thruster:smallentity:ship-part:thruster:small entity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:hull:triangle #entity:ship-part:weapon:mass-driverentity:ship-part:hull:square #entity:ship-part:weapon:mass-driverentity:ship-part:thruster:smallentity:ship-part:thruster:small  hexagon   entity:ship-part:hull:square entity:ship-part:hull:triangle    entity:ship-part:hull:triangle entity:ship-part:hull:square  entity:ship-part:hull:triangle  entity:ship-part:hull:hexagon  entity:ship-part:hull:square  entity:ship-part:hull:hexagon    entity:ship-part:hull:triangle entity:ship-part:hull:square  entity:ship-part:hull:triangle  entity:ship-part:hull:hexagon  entity:ship-part:hull:square  entity:ship-part:hull:hexagon    entity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:small                  entity:ship-part:hull:triangle entity:ship-part:hull:hexagon   entity:ship-part:hull:square  entity:ship-part:hull:hexagon   entity:ship-part:hull:square entity:ship-part:thruster:small entity:ship-part:hull:triangle   entity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:small       entity:ship-part:hull:square  entity:ship-part:hull:triangle  entity:ship-part:hull:square      mallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:small  entity:ship-part:hull:triangle entity:ship-part:hull:triangle entity:ship-part:hull:triangle   entity:ship-part:hull:triangle  entity:ship-part:hull:triangle entity:ship-part:hull:square  entity:ship-part:hull:triangle  entity:ship-part:hull:square         entity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:small#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driverentity:ship-part:hull:square #entity:ship-part:weapon:mass-driverentity:ship-part:hull:triangle #entity:ship-part:weapon:mass-driverentity:ship-part:hull:triangle entity:ship-part:hull:triangle #entity:ship-part:weapon:mass-driverentity:ship-part:hull:triangle entity:ship-part:hull:triangle #entity:ship-part:weapon:mass-driverentity:ship-part:hull:triangle entity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:hull:triangle entity:ship-part:thruster:smallentity:ship-part:hull:hexagon entity:ship-part:thruster:smallentity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:hull:hexagon  entity:ship-part:thruster:smallentity:ship-part:hull:hexagon entity:ship-part:hull:triangle  entity:ship-part:hull:triangle entity:ship-part:hull:triangle entity:ship-part:hull:triangle  entity:ship-part:hull:square  entity:ship-part:hull:triangle     entity:ship-part:hull:triangle    entity:ship-part:hull:square entity:ship-part:hull:square  entity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:hull:triangle entity:ship-part:thruster:smallentity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:hull:triangle entity:ship-part:hull:hexagon entity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:hull:hexagon entity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:small  entity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:hull:square entity:ship-part:thruster:small entity:ship-part:thruster:smallentity:ship-part:thruster:small  entity:ship-part:hull:triangle entity:ship-part:hull:triangle entity:ship-part:hull:triangle   entity:ship-part:hull:triangle  entity:ship-part:hull:triangle entity:ship-part:hull:square  entity:ship-part:hull:triangle  entity:ship-part:hull:square  entity:ship-part:hull:triangle entity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:hull:triangle entity:ship-part:thruster:smallentity:ship-part:hull:hexagon entity:ship-part:thruster:smallentity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:hull:hexagon  entity:ship-part:hull:square  entity:ship-part:hull:square entity:ship-part:hull:triangle entity:ship-part:thruster:smallentity:ship-part:hull:hexagon entity:ship-part:thruster:small entity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:hull:hexagon entity:ship-part:thruster:small entity:ship-part:hull:square entity:ship-part:hull:triangle entity:ship-part:thruster:small  #entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver  #entity:ship-part:weapon:mass-driver #entity:ship-part:weapon:mass-driverentity:ship-part:hull:triangle entity:ship-part:hull:hexagon  #entity:ship-part:weapon:mass-driverentity:ship-part:hull:square  entity:ship-part:hull:hexagon  #entity:ship-part:weapon:mass-driverentity:ship-part:hull:square #entity:ship-part:weapon:mass-driverentity:ship-part:hull:square  entity:ship-part:hull:square entity:ship-part:hull:triangle entity:ship-part:thruster:smallentity:ship-part:hull:hexagon entity:ship-part:thruster:small entity:ship-part:hull:square entity:ship-part:thruster:smallentity:ship-part:hull:hexagon entity:ship-part:thruster:small entity:ship-part:hull:square entity:ship-part:hull:triangle entity:ship-part:thruster:small  #entity:ship-part:weapon:mass-driver#entity:ship-part:weapon:mass-driver  #entity:ship-part:weapon:mass-driver #entity:ship-part:weapon:mass-driverentity:ship-part:hull:triangle entity:ship-part:hull:hexagon  #entity:ship-part:weapon:mass-driverentity:ship-part:hull:square  entity:ship-part:hull:hexagon  #entity:ship-part:weapon:mass-driverentity:ship-part:hull:square #entity:ship-part:weapon:mass-driver entity:ship-part:hull:triangle  entity:ship-part:thruster:small entity:ship-part:thruster:smallentity:ship-part:thruster:small entity:ship-part:thruster:smallentity:ship-part:thruster:small entity:ship-part:hull:triangle  entity:ship-part:thruster:small entity:ship-part:thruster:smallentity:ship-part:thruster:small entity:ship-part:thruster:smallentity:ship-part:thruster:small entity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:small    entity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:smallentity:ship-part:thruster:small    entity:ship-part:hull:square #entity:ship-part:weapon:mass-driverentity:ship-part:hull:triangle #entity:ship-part:weapon:mass-driver   entity:ship-part:thruster:smallentity:ship-part:thruster:small