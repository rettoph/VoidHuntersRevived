ship-part:chassis:mosquitoship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:small ship-part:hull:pentagon   ship-part:weapon:mass-driver ship-part:weapon:mass-drivership-part:hull:pentagon  ship-part:weapon:mass-driver   hull:pentagon ship-part:thruster:smallship-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:hull:pentagon ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:smallship-part:thruster:small lship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:smallship-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-driver  ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:pentagon ship-part:weapon:mass-drivership-part:square  ship-part:beam:horizontalship-part:thruster:small   ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:square ship-part:thruster:smallship-part:beam:horizontal   ship-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:smallship-part:thruster:small ship-part:thruster:smallship-part:thruster:small pon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:smallship-part:thruster:smallship-part:thruster:small :pentagonship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:weapon:mass-drivership-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:thruster:smallship-part:pentagonship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:thruster:smallship-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:smallship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:squareship-part:weapon:mass-drivership-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:squareship-part:weapon:mass-drivership-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-driver ship-part:thruster:smallship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:pentagonship-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:thruster:smallship-part:pentagonship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:thruster:smallship-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:smallship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:squareship-part:weapon:mass-drivership-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:squareship-part:weapon:mass-drivership-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:thruster:smallship-part:pentagonship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:thruster:smallship-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:smallship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:squareship-part:weapon:mass-drivership-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:squareship-part:weapon:mass-drivership-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-driver ship-part:thruster:small