ship-part:hull:hexagonship-part:hull:pentagon   ship-part:hull:square  ship-part:hull:hexagon  ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:hull:pentagon ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:hull:square ship-part:weapon:mass-driver      ship-part:hull:pentagon   ship-part:hull:square  ship-part:hull:hexagon  ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:hull:pentagon ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:hull:square ship-part:weapon:mass-driver      ship-part:hull:pentagon   ship-part:hull:square  ship-part:hull:hexagon  ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:hull:pentagon ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:hull:square ship-part:weapon:mass-driver      ship-part:hull:pentagon   ship-part:hull:square  ship-part:hull:hexagon  ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:hull:pentagon ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:hull:square ship-part:weapon:mass-driver      ship-part:hull:pentagon   ship-part:hull:square  ship-part:hull:hexagon  ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:hull:pentagon ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:hull:square ship-part:weapon:mass-driver      ship-part:hull:pentagon   ship-part:hull:square  ship-part:hull:hexagon  ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:hull:pentagon ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:hull:square ship-part:weapon:mass-driver      rt:thruster:small ship-part:thruster:smallship-part:thruster:smallship-part:hull:square  ship-part:hull:pentagon  ship-part:hull:pentagon  ship-part:hull:pentagon ship-part:thruster:smallship-part:hull:square ship-part:thruster:small ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:small ship-part:thruster:smallship-part:thruster:smallhruster:smallship-part:thruster:smallss-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:square  ship-part:beam:horizontalship-part:thruster:small ship-part:thruster:small ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-driver  ship-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-driver  ship-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-drivership-part:pentagon ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:smallship-part:thruster:small  ship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:weapon:mass-driver     ship-part:weapon:mass-driver  mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:thruster:smallship-part:pentagonship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:squareship-part:weapon:mass-drivership-part:pentagonship-part:thruster:smallship-part:pentagonship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:thruster:smallship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:squareship-part:weapon:mass-drivership-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:squareship-part:weapon:mass-drivership-part:thruster:smallship-part:pentagonship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:weapon:mass-drivership-part:weapon:mass-drivership-part:squareship-part:weapon:mass-driver ship-part:thruster:small ship-part:thruster:small