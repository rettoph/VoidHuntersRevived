 Unnamed Shipvhr:chassis:fightervhr:weapon:mass-driver:tinyvhr:thruster:tinyvhr:thruster:tinyvhr:thruster:tinyvhr:thruster:tiny