ship-part:chassis:mosquitoship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:smallship-part:thruster:small ship-part:pentagon  ship-part:weapon:mass-driver ship-part:weapon:mass-drivership-part:pentagon ship-part:weapon:mass-driver   smallship-part:thruster:smallship-part:weapon:mass-driver ship-part:weapon:mass-drivership-part:pentagon ship-part:weapon:mass-drivership-part:thruster:smallship-part:thruster:small 