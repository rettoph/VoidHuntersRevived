 Unnamed Shipvhr:chassis:waspvhr:hull:pentagonvhr:weapon:mass-driver vhr:thruster:smallvhr:thruster:smallvhr:thruster:smallvhr:weapon:mass-drivervhr:thruster:small        vhr:thruster:smallvhr:weapon:mass-drivervhr:thruster:small  vhr:thruster:small  vhr:weapon:mass-drivervhr:hull:pentagonvhr:thruster:smallvhr:thruster:smallvhr:weapon:mass-driver     